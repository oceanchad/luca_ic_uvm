`include "param_def.v"

