module factory_override;
    import uvm_pkg::;
    
endmodule