`include "param_def.v"

package mcdf_pkg;
    import chnl_pkg::*;
    import reg_pkg::*;
    import arb_pkg::*;
    import fmt_pkg::*;
    import rpt_pkg::*;

    
endpackage