`ifndef APB_SVH
`define APB_SVH

`include "apb_transfer.svh"
`include "apb_config.sv"

`include "apb_master_driver.svh"
`include "apb_master_monitor.svh"
`include "apb_master_sequencer.svh"
`include "apb_master_agent.svh"

